//`infdef APB_PKG
//`define APB_PKG
 package apb_pkg;
   event e1; 
   `include "/home/dvft0901/apb_sv_project/env/apb_transaction.sv"
   `include "/home/dvft0901/apb_sv_project/env/apb_generator.sv"   
   `include "/home/dvft0901/apb_sv_project/env/apb_driver.sv"
   `include "/home/dvft0901/apb_sv_project/env/apb_monitor.sv"
   `include "/home/dvft0901/apb_sv_project/env/apb_predictor.sv" 
   `include "/home/dvft0901/apb_sv_project/env/apb_scoreboard.sv"   
   `include "/home/dvft0901/apb_sv_project/env/apb_enviroment.sv"   
   `include "/home/dvft0901/apb_sv_project/test/apb_test.sv"

endpackage 
