//`infdef APB_PKG
//`define APB_PKG
 package apb_pkg;
   event e1; 
   `include "apb_transaction.sv"
   `include "apb_generator.sv"   
   `include "apb_driver.sv"
   `include "apb_monitor.sv"
   `include "apb_predictor.sv" 
   `include "apb_scoreboard.sv"   
   `include "apb_enviroment.sv"   
   `include "apb_test.sv"

endpackage 
